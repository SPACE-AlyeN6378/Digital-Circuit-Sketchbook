library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


-- ============================================================================
entity {entity_name} is
    port (
        {port_declarations}
    );
end entity {entity_name};
-- ============================================================================

architecture {architecture_name} of {entity_name} is
    {signal_declarations}
    
begin
    {gate_operations}

end {architecture_name};
    
